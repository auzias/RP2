library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY test_bench_half_adder IS
END test_bench_half_adder;