architecture ha of halfAdder is

begin
	S <= A xor B;
	Cy <= A and B;
end ha;
