library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity test_bench_mux is
end test_bench_mux;